Author: Manish Singhal
Date: 2nd Mar 15


class producer extends uvm_component;
// $display
endclass: producer


class consumer extends uvm_component;

endclass: consumer

class env extends uvm_env;

endclass: env
